LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ROM IS
	PORT(
		entrada : IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		saida	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END ROM;

ARCHITECTURE arch OF ROM IS
BEGIN
	WITH entrada SELECT
	--  saida <=    "DADO_MEM" WHEN "ADDR_MEM",
		saida <= 	"00101010" WHEN "00000000",
					"01111111" WHEN "00000001",
					"01010111" WHEN "00000010",
					"00101111" WHEN "00000011",
					"01110101" WHEN "00000100",
					"01111101" WHEN "00000101",
					"01111001" WHEN "00000110",
					"00000000" WHEN OTHERS;
END arch; 